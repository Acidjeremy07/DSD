library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SRLATCH is
	port (	S	:	IN	STD_LOGIC;
			R	:	IN	STD_LOGIC;
			XA	:	OUT	STD_LOGIC;
			XB	:	OUT STD_LOGIC;
			MXA	:	IN	STD_LOGIC;
			MXB	:	IN	STD_LOGIC;
			MS	:	IN	STD_LOGIC);

ATTRIBUTE PIN_NUMBERS OF SRLATCH: ENTITY IS
	" S:2 R:3 MS:4 MXA:5 MXB:6 "
	& " XA:14 XB:15 ";

END SRLATCH;


ARCHITECTURE FUNCION OF SRLATCH IS 
	SIGNAL	notQ	:	STD_LOGIC;
	SIGNAL	Q		:	STD_LOGIC;
	SIGNAL	MUXOUT	:	STD_LOGIC;
	BEGIN

		Q<= R nor notQ;
		notQ<= S nor notQ;

		MUXOUT<= (NOT MS AND MXA) OR (MS AND MXB);
	
		XA<= Q AND MUXOUT;
		XB<= notQ AND MUXOUT;

END FUNCION;

		
